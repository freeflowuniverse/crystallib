module tfgrid

pub struct KeyValue {
pub mut:
 	key string
	value string
}
