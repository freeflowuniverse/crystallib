module bizmodel

