module data
