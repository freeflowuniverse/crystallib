module taiga

import json

struct Story {
pub mut:
	description            string
	id                     int
	is_private             bool
	tags                   []string
	project                int
	project_extra_info     ProjectInfo
	status                 int
	status_extra_info      StatusInfo
	assigned_to            int
	assigned_to_extra_info UserInfo
	owner                  int
	owner_extra_info       UserInfo
	created_date           string
	modified_date          string
	finish_date            string
	subject                string
	is_closed              bool
	is_blocked             bool
	blocked_note           string
	ref                    int
	client_requirement     bool
	team_requirement       bool
	tasks                  []Task
}

struct NewStory {
pub mut:
	subject string
	project int
}

pub fn (mut h TaigaConnection) stories() ?[]Story {
	data := h.get_json_str('stories', '', true) ?
	return json.decode([]Story, data) or {}
}

pub fn (mut h TaigaConnection) story_create(subject string, project_id int) ?Story {
	h.cache_drop()? //to make sure all is consistent
	story := NewStory{
		subject: subject
		project: project_id
	}
	postdata := json.encode_pretty(story)
	response := h.post_json_str('stories', postdata, true, true) ?
	mut result := json.decode(Story, response) ?
	return result
}

pub fn (mut h TaigaConnection) story_get(id int) ?Story {
	// TODO: Check Cache first (Mohammed Essam)
	response := h.get_json_str('stories/$id', "", true) ?
	mut result := json.decode(Story, response) ?
	return result
}
