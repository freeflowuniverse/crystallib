module analytics

pub enum Event {
	custom
	http_request
}
