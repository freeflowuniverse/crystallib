module coinmarketcap
module gittools

import os

fn test_1() {
	
	panic("sss")

}