module tailwind


[heap]
pub struct TailwindFactory {
pub mut:
}

pub fn new() TailwindFactory {
	mut twf:=TailwindFactory{}
	return twf
}
