module encoderhero

import time
