module smartid

import freeflowuniverse.crystallib.redisclient


fn test_load() {
	defer {
		cleanup(mut redis) or { panic(err) }
	}

	t:='
	
'
	//TODO: sid_empty_replace
	
}
