module testactor

pub struct BaseObject {
	text string @[index]
	number int
}

