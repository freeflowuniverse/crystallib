module syncthing

fn (mut a App) deploy() ! {
}
