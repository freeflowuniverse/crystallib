module generic

// import freeflowuniverse.crystallib.ui.console
// import freeflowuniverse.crystallib.ui.telegram { UITelegram }
import freeflowuniverse.crystallib.ui.uimodel

// ...
// ```
// args:
// TODO
// }
// ```
pub fn (mut c UserInterface) pay(args uimodel.PayArgs) ! {
	// match mut c.channel {
	// 	UIConsole { return c.channel.editor(args)! }
	// 	else { panic("can't find channel") }
	// }
}
