module circles

// pub struct BusinessModel {
// 	employees
// }
