module twinsafe

//TODO: create 2 tables, one for othertwin, one for mytwin