module zos

pub struct ZOSClient {
}
