module template

import freeflowuniverse.crystallib.ui.uimodel { QuestionArgs }

pub fn (mut c UIExample) ask_date(args QuestionArgs) string {
	panic('implement')
}

pub fn (mut c UIExample) ask_time(args QuestionArgs) string {
	panic('implement')
}
