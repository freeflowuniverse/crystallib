module builder

[heap]
pub struct NodesFactory {
pub mut:
	nodes map[string]&Node
}
