module planner

import texttools

// texttools.text_to_params()?
