module publisher2

import freeflowuniverse.crystallib.publisher2

fn do() ? {

}

fn main() {
	do() or { panic(err) }
}
