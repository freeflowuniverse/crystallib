module syncthing

const name="syncthing"
