module data

//Data object for User
pub struct User {
pub mut:
	id          int
	name        string
	description string
	tags		[]string
	remarks		[]int
}