module people

import freeflowuniverse.crystallib.baobab.models.system
import json

fn test_1() {
	mut p := person_new()?
	// p.start_date.now()

	// println(p)

	// panic('s')
}
