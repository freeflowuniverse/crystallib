module project

pub enum State {
	new
	active
	blocked
	done
	verified
}

pub enum Priority {
	low
	normal
	urgnet
}
