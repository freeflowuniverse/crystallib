module webserver
