module backoffice

