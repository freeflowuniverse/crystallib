module calc
