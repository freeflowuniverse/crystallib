module encoder


fn test_encode() {}


fn test_decode() {}