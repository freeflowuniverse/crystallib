module budget

//! This seems redundant, we can just use the budget_item_person.v file
