module installers

// following functions are set of utilities to make our life easy, use vlang as constructs (not the builder)
