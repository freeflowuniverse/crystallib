module grid

fn test_vm_deploy() ! {
	deployer := new_deployer('license carry boss sand squeeze forum wide try reform embrace chimney mimic brass wreck wing dove tiger admit jelly quit water twist face pull')!
	deployer.vm_deploy(
		name: 'test_vm'
		deployment_name: 'test_deployment'
	)
}