module play

pub struct Base {
pub mut:
	session ?&Session @[skip; str: skip]
	name    string
}

pub fn (mut self Base) session() !&Session {
	mut session := self.session or {
		mut s := session_new()!
		self.session = s
		s
	}

	return session
}

pub fn (mut self Base) context() !&Context {
	mut session := self.session()!
	return &session.context
}
