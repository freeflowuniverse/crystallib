module gittools

import os
import freeflowuniverse.crystallib.osal
import freeflowuniverse.crystallib.ui.console
import freeflowuniverse.crystallib.core.pathlib
import freeflowuniverse.crystallib.core.base
import freeflowuniverse.crystallib.develop.vscode
import freeflowuniverse.crystallib.develop.sourcetree

@[heap]
pub struct GitRepo {
	id int
pub mut:
	gs   &GitStructure @[skip; str: skip]
	addr &GitAddr
	status &GitRepoStatus
	path pathlib.Path
}


pub fn (repo GitRepo) key() string {
	return repo.addr.key()
}

fn ( repo GitRepo) cache_key() string {
	return '${gitstructure_key(repo.gs.coderoot.path)}:${repo.addr.provider}:${repo.addr.account}:${repo.addr.name}'
}

// remove cache
pub fn (repo GitRepo) cache_delete() ! {
	mut c := base.context()!
	mut redis := c.redis()!	
	redis.del(repo.cache_key())!
}


pub fn (mut repo GitRepo) load() !GitRepoStatus {
	repo.path.check() // could be that path changed
	if !repo.path.exists() {
		return error("cannot load from path, doesn't exist for '${repo.path.path}'")
	}

	// TODO: fix
	// mut c := base.context()!
	// mut redis := c.redis()!
	// mut isvalid := redis.get(repo.addr.cache_key_status() + '_') or { '' }
	// if isvalid != '' {
	// 	return repo.status()!
	// }
	mut st := repo_load(mut repo.addr, repo.path.path)!
	repo.status_set(st)!

	p2 := repo.addr.path()!
	if p2.path != repo.path.path {
		return error("path conflict, doesn't exist for '${p2.path}' and '${repo.path.path}'")
	}
	// console.print_header(' status:\n${st}')
	// redis.set(repo.addr.cache_key_status() + '_', '1')!
	// redis.expire(repo.addr.cache_key_status() + '_', 5)! // 5 seconds, to not have these double gets
	return st
}

pub fn (mut repo GitRepo) need_pull() !bool {
	s := repo.status()!
	return s.need_pull
}

// relative path inside the gitstructure, pointing to the repo
pub fn (repo GitRepo) path_relative() string {
	return repo.path.path_relative(repo.gs.coderoot.path) or { panic('couldnt get relative path') } // TODO: check if works well
}

// pulls remote content in, will reset changes
pub fn (mut repo GitRepo) pull_reset(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	repo.remove_changes(args)!
	repo.pull(args)!
}

@[params]
pub struct ActionArgs {
pub mut:
	reload bool = true
	msg    string // only relevant for commit
	branch string
	tag string
	recursive bool
}

// commit the changes, message is needed, pull from remote, push to remote
pub fn (mut repo GitRepo) commit_pull_push(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	repo.commit(args)!
	repo.pull(args)!
	repo.push(args)!
}

// commit the changes, message is needed, pull from remote
pub fn (mut repo GitRepo) commit_pull(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	repo.commit(args)!
	repo.pull(args)!
}

// pulls remote content in, will fail if there are local changes
pub fn (mut repo GitRepo) pull(args_ ActionArgs) ! {
	$if debug {
		console.print_debug('  pull: ${repo.url_get(true)} (branch: ${args_.branch})')
	}
	// repo.ssh_key_load()!
	// defer {
	// 	repo.ssh_key_forget() or { panic("bug") }
	// }

	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}

	
	if args.branch != '' {
		//console.print_debug(" - branch detected: '${repo.addr.branch}'")
		if args.branch != repo.addr.branch  {
			console.print_header(' branch pull ${repo.addr.branch} -> ${args.branch} for ${repo.addr.remote_url}')
			repo.branch_switch(args.branch)!
		}
	}

	// } else {
	// 	print_backtrace()
	// 	return error('branch should have been known for ${repo.addr.remote_url}')

	// st := repo.status()!
	// if st.need_commit {
	// 	return error('Cannot pull repo: ${repo.path.path}, a commit is needed.\n${st}')
	// }
	// pull can't see the status
	cmd2 := 'cd ${repo.path.path} && git pull'
	osal.execute_silent(cmd2) or {
		console.print_debug(' GIT PULL FAILED: ${cmd2}')
		return error('Cannot pull repo: ${repo.path}. Error was ${err}')
	}

	if args.tag != '' {
		console.print_header("tag pull: '${args.tag}' for ${repo.addr.remote_url} ")
		cmd := 'cd ${repo.path.path} && git checkout ${args.tag}'
		osal.execute_silent(cmd) or {
			return error('Cannot pull tag ${args.tag} for  repo: ${repo.path.path}. \nError was ${err}')
		}
	}

	if args.recursive{
		cmd3:="cd ${repo.path.path} && git submodule update --init --recursive"
		osal.execute_silent(cmd3) or {
			console.print_debug(' GIT RECURSIVE PULL FAILED: ${cmd3}')
			return error('Cannot pull repo: ${repo.path}. Error was ${err}')
		}		
	}
	repo.load()!

	// repo.ssh_key_forget()!
}

// pub fn (mut repo GitRepo) rev() !string {
// 	// $if debug {
// 	// 	console.print_debug('   - REV: ${repo.url_get(true)}')
// 	// }
// 	cmd2 := 'cd ${repo.path.path} && git rev-parse HEAD'
// 	res := osal.execute_silent(cmd2) or {
// 		console.print_debug(' GIT REV FAILED: ${cmd2}')
// 		return error('Cannot rev repo: ${repo.path}. Error was ${err}')
// 	}
// 	return res.trim_space()
// }

pub fn (mut repo GitRepo) commit(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	st := repo.status()!
	if st.need_commit {
		if args.msg == '' {
			return error('Cannot commit, message is empty for ${repo}')
		}
		cmd := "
		cd ${repo.path.path}
		set +e
		git add . -A
		git commit -m \"${args.msg}\"
		echo "
		osal.execute_silent(cmd) or {
			return error('Cannot commit repo: ${repo.path.path}. Error was ${err}')
		}
	} else {
		console.print_debug('     > no change')
	}
	repo.load()!
}

// remove all changes of the repo, be careful
pub fn (mut repo GitRepo) remove_changes(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	st := repo.status()!
	if st.need_commit {
		console.print_header(' remove change ${repo.path.path}')
		cmd := '
		cd ${repo.path.path}
		rm -f .git/index
		#git fetch --all
		git reset HEAD --hard
		git clean -xfd		
		git checkout . -f
		echo ""
		'
		res := osal.exec(cmd: cmd, raise_error: false)!
		console.print_debug(cmd)
		// console.print_debug(res)
		if res.exit_code > 0 {
			console.print_header(' could not remove changes, will re-clone ${repo.path.path}')
			repo.path.delete()! // remove path, this will re-clone the full thing
			repo.load_from_url()!
		}
	}
	repo.load()!
}

pub fn (mut repo GitRepo) push(args_ ActionArgs) ! {
	mut args := args_
	if args.reload {
		repo.load()!
		args.reload = false
	}
	$if debug {
		console.print_debug('   - PUSH: ${repo.url_get(true)} on ${repo.path.path}')
	}
	// repo.ssh_key_load()!
	// defer {
	// 	repo.ssh_key_forget() or { panic(err) }
	// }
	st := repo.status()!
	if st.need_push {
		console.print_debug('    - PUSH THE CHANGES')
		cmd := 'cd ${repo.path.path} && git push'
		osal.execute_silent(cmd) or {
			return error('Cannot push repo: ${repo.path.path}. Error was ${err}')
		}
	}
	repo.load()!
	// repo.ssh_key_forget()!
}

pub fn (mut repo GitRepo) branch_switch(branchname string) ! {
	if repo.gs.config.multibranch {
		return error('cannot do a branch switch if we are using multibranch strategy.')
	}
	repo.load()!
	st := repo.status()!
	if st.need_commit || st.need_push {
		return error('Cannot branch switch repo: ${repo.path.path} because there are changes in the dir.')
	}
	// Fetch repo before checkout, in case a new branch added.
	repo.fetch_all()!
	cmd := 'cd ${repo.path.path} && git checkout ${branchname}'
	osal.execute_silent(cmd) or {
		// console.print_debug('GIT CHECKOUT FAILED: $cmd_checkout')
		return error('Cannot branch switch repo: ${repo.path.path}. Error was ${err} \n cmd: ${cmd}')
	}
	// console.print_debug(cmd)
	repo.pull(reload: true)!
}

pub fn (mut repo GitRepo) fetch_all() ! {
	// repo.ssh_key_load()!
	// defer {
	// 	repo.ssh_key_forget() or { panic(err) }
	// }
	cmd := 'cd ${repo.path.path} && git fetch --all'
	osal.execute_silent(cmd) or {
		// console.print_debug('GIT FETCH FAILED: $cmd_checkout')
		return error('Cannot fetch repo: ${repo.path.path}. Error was ${err} \n cmd: ${cmd}')
	}
	repo.load()!
	// repo.ssh_key_forget()!
}

// deletes git repository
pub fn (mut repo GitRepo) delete() ! {
	$if debug {
		console.print_debug('   - DELETE: ${repo.url_get(true)}')
	}
	if !os.exists(repo.path.path) {
		return
	} else {
		panic('implement')
	}
	repo.cache_delete()!
}

//////////////////////////KEY MGMT
//////////////////////////////////

// set the key (private ssh key)
pub fn (repo GitRepo) ssh_key_set(key string) ! {
	mut p := pathlib.get_file(path: repo.ssh_key_path(), create: true)!
	p.write(key)!
}

fn (repo GitRepo) ssh_key_path() string {
	return '${os.home_dir()}/.ssh/${repo.key()}'
}

//////////////////////////EDIT CODE MGMT
//////////////////////////////////

// open sourcetree for the git repo
pub fn (repo GitRepo) sourcetree() ! {
	sourcetree.open(path: repo.path.path)!
}

// open visual studio code for repo
pub fn (repo GitRepo) vscode() ! {
	vscode.open(path: repo.path.path)!
}
