module processmanager

import freeflowuniverse.crystallib.osal

pub struct ProcessManager {
	// pub mut:
}

pub fn new() !ProcessManager {
	mut pm := ProcessManager{}
}
