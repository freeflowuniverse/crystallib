module zola

fn test_section_export() {
	section := Section{}
	section.export('test')!
<<<<<<< HEAD
<<<<<<< HEAD
}
=======
}
>>>>>>> e61681d (example fix wip)
=======
}
>>>>>>> 2007ff6 (fix sections processing)
