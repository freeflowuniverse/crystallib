module books

[heap]
pub struct Config {
pub mut: // pointer to site
	heal bool = true
	dest string = "/tmp/mdbooks"
	mdbook_template_path string 
}
