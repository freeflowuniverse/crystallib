module openrpc

// pub struct 