module installers

import freeflowuniverse.crystallib.core.pathlib
import freeflowuniverse.crystallib.osal.gittools
