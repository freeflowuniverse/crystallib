module base

__global (
	contexts        map[u32]&Context
	context_current u32
)
