module blockchain

// import freeflowuniverse.crystallib.data.actionsparser

pub struct Controller {
}

pub fn new() !Controller {
	mut c := Controller{}
	return c
}
