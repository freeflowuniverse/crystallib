module petstore_client

// a pet struct that represents a pet
struct Pet {
	name string // name of the pet
	tag  string // a tag of the pet, helps finding pet
	id   int    // unique indentifier
}
