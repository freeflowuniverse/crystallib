module books

[heap]
struct MDBookInstance {
mut:
	name string
}
