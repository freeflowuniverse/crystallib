module tasklets

//@for domainname,domain in tm.domains
//@for actorname,actor in domain.actors
// import domain_@{domainname}.actor_@{actorname}
//@end
//@end

// fn (mut tm &TaskletManager) action_reboot(mut job &actionrunner.ActionJob)!bool{
