module vbuilder

const name = 'vbuilder'
