module servers
