module currency

pub struct Currency {
pub mut:
	name   string
	usdval f64
}
