module builder

fn test_nodedb() {
	// TODO URGENT create tests for nodedb
}

fn test_nodedone() {
	// TODO URGENT create tests for nodedone
}
