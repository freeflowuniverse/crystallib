module jobs

import freeflowuniverse.crystallib.data.paramsparser
import time
