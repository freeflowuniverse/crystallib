module griddriver

pub struct Client {
pub:
	mnemonic  string
	substrate string
	relay     string
}

// TODO: add the rest of griddriver functionalities
