module model

[root ; inherit:'base']
pub struct Group {
pub mut:
	users	[]u32
}

