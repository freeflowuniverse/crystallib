module lima

cmd = 'limactl create default --cpus 16 --memory 4 --containerd system'
