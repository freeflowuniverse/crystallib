module threefold
