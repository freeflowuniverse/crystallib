module jsonschema

fn test_define() {
	mut schema := Schema{}
	// schema.define()
}