module components

import db.sqlite
import nedpals.vex.ctx

fn get_db(req &ctx.Req) ?&sqlite.DB {
	raw_db := req.ctx.value('db')?
	if raw_db is sqlite.DB {
		return raw_db
	}
	return none
}
