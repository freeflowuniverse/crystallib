module publishermod

import texttools
import os

// the factory, get your tools here
// use path="" if you want to go from os.home_dir()/code/
// will find all wiki's
pub fn new(path string) ?Publisher {
	mut publisher := Publisher{}
	publisher.gitlevel = 0
	publisher.replacer.site = texttools.regex_instructions_new() or { panic(err) }
	publisher.replacer.file = texttools.regex_instructions_new() or { panic(err) }
	publisher.replacer.word = texttools.regex_instructions_new() or { panic(err) }
	publisher.find_sites(path.replace('~', os.home_dir())) ?

	return publisher
}

// check all pages, try to find errors
pub fn (mut publisher Publisher) check() {
	for mut site in publisher.sites {
		site.load(mut publisher)
	}
	for mut site in publisher.sites {
		site.process(mut publisher)
	}
	publisher.defs_pages_init()
}

// returns the found locations for the sites, will return [[name,path]]
pub fn (mut publisher Publisher) site_locations_get() [][]string {
	mut res := [][]string{}
	for site in publisher.sites {
		res << [site.name, site.path]
	}
	return res
}
