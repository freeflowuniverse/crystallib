module jobs

import freeflowuniverse.crystallib.params
import time
