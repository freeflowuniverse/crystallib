module milvus
