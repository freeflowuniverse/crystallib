module publisher2


// install mdbook will return true if it was already installed
pub fn get() ?Publisher {
	mut p := Publisher{
	}
	return p
}