module tools
