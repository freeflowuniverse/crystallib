module main



fn main() {

}
