module vdc

pub struct DISK {
pub mut:
	name        string
	description string
}
