module main

import freeflowuniverse.crystallib.verasure

fn main() {

	verasure.test()
	// mut e := verasure.new(16, 4)
	// shards := e.encode('Lorem ipsum dolor sit amet, consectetur adipiscing elit. Integer consectetur accumsan augue, at pharetra'.bytes())
	// println(shards)

	// data := e.decode(shards)
	// println(data.len)
	// println(data.bytestr())


}
