module vbuilder



fn (mut a App) deploy() !{

	

}