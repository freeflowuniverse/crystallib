module calc

