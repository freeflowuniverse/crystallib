module stellar


