module gittools

import freeflowuniverse.crystallib.pathlib

