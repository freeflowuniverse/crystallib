module usermanager



pub struct Contact {
pub mut:

	name string 
}

