module installers

// import freeflowuniverse.crystallib.core.pathlib
// import freeflowuniverse.crystallib.develop.gittools

@[params]
pub struct UploadArgs {
pub mut:
	cmdname string
	source  string
	reset   bool
}

pub fn upload(args_ UploadArgs) ! {
	mut args := args_
	panic('to implement')
}
