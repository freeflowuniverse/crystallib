module blockchain

// import freeflowuniverse.crystallib.data.actionparser

pub struct Controller {
}

pub fn new() !Controller {
	mut c := Controller{}
	return c
}
