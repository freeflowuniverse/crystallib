module analytics

// import db.sqlite

// @[params]
// pub struct DBBackendConfig {
// 	db_path string = 'analytics.sqlite'
// }

// // factory for
// pub fn new_backend(config DBBackendConfig) !DBBackend {
// 	db := sqlite.connect(config.db_path) or { panic(err) }

// 	sql db {
// 		create table Log
// 	} or { panic(err) }

// 	return DBBackend{
// 		db: db
// 	}
// }
