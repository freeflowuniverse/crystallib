module params


pub fn (mut result Params) str()string {
	//TODO: walk over params fill in a serialized string
	//TODO: Jonathan
	return ""
}
