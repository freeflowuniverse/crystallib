module liquid
module gittools

import os

fn test_1() {

	// key = "92be9b29-7f6c-48e4-9ef2-d6aa0550f620"

	mut c := new({secret:key})

	//need to fetch USD/TFT price
	//see how we did for taiga how to use the connection



	panic("sss")

}