module backoffice
