module data

//Data object for Circle
pub struct Circle {
pub mut:
	id          int
	name        string
	description string
	tags		[]string
	remarks		[]int
}