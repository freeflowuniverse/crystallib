module resp

import io

// fn print_val_to_check(s string) {
// 	println(s.replace('\n', '\\\\n').replace('\r', '\\\\r'))
// }
