module pathlib

import os

// gets Path object, will check if it exists, is dir_file, ...
pub fn get(path_ string) Path {
	mut path := path_
	if path.contains('~') {
		path = path.replace('~', os.home_dir())
	}
	if path.contains('file://') {
		path = path.trim_string_left('file://')
	}
	mut p2 := Path{
		path: path
	}
	p2.check()
	if p2.path.contains('..') {
		p2.path = p2.absolute()
	}
	return p2
}

pub fn get_no_check(path string) Path {
	mut p2 := Path{
		path: path
	}
	return p2
}

[params]
pub struct GetArgs{
pub mut:
	path string
	create bool
	check bool = true //means will check the dir or file exists
	empty bool //will empty the dir or the file
}

// get a directory, or needs to be created
// if the dir doesn't exist and is not created, then there will be an error
pub fn get_dir(args_ GetArgs) !Path {
	mut args:=args_
	if args.empty{
		args.create=true
	}		
	if args.create{
		args.check=true
	}
	mut p2 := get(args.path)
	if args.check{
		// p2.check()
		p2.absolute()
		if p2.exist == .no {
			os.mkdir_all(p2.absolute()) or { return error('cannot create path ${p2}') } // Make sure that all the needed paths created		
			p2.check()
		}
		if !p2.is_dir() {
			return error('Path ${args.path} is not a dir.')
		}
		if args.empty{
			p2.empty()!
		}
	}
	return p2
}

pub fn get_file(args_ GetArgs) !Path {
	mut args:=args_
	if args.empty{
		args.create=true
	}		
	if args.create{
		args.check=true
	}
	mut p2 := get(args.path)
	if args.check{
		// p2.check()
		if args.create{
			parent_ := p2.parent()!
			if parent_.exist == .no {
				os.mkdir_all(parent_.path) or { return error('cannot create path:${args.path}') }
			}
			if p2.exist == .no ||  args.empty{
				os.write_file(args.path, '') or { return error('cannot create empty file:${args.path}') }
				p2.check()
			}
		}
		if !p2.is_file() {
			return error('Path ${args.path} is not a file.')
		}		
	}
	return p2
}
