module jobs

