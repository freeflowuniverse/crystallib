module peertube

import freeflowuniverse.crystallib.installers.base
import freeflowuniverse.crystallib.tools.tmux
import freeflowuniverse.crystallib.osal
import freeflowuniverse.crystallib.core.pathlib
import freeflowuniverse.crystallib.core.texttools
import os

[params]
pub struct InstallArgs {
pub mut:
	reset bool
}

// TODO: make installer for peertube

// install peertube will return true if it was already installed
pub fn install(args InstallArgs) ! {
	// make sure we install base on the node
	base.install()!

	if args.reset == false && osal.done_exists('install_peertube') {
		return
	}

	// install peertube if it was already done will return true
	println(' - package_install install peertube')

	if osal.platform() != .ubuntu {
		return error('only support ubuntu for now')
	}
	// mut dest := osal.download(
	// 	url: 'https://github.com/peertubeserver/peertube/releases/download/v2.7.4/peertube_2.7.4_linux_amd64.tar.gz'
	// 	minsize_kb: 10000
	// 	reset: true
	// 	expand_dir: '/tmp/peertubeserver'
	// )!

	// mut peertubefile := dest.file_get('peertube')! // file in the dest
	// peertubefile.copy('/usr/local/bin')!
	// peertubefile.chmod(0o770)! // includes read & write & execute

	// osal.done_set('install_peertube', 'OK')!
	return
}

[params]
pub struct WebConfig {
pub mut:
	path   string = '/var/www'
	domain string = ''
}

// configure peertube as default webserver & start
// node, path, domain
// path e.g. /var/www
// domain e.g. www.myserver.com
pub fn configure_examples(config WebConfig) ! {
	mut config_file := $tmpl('templates/peertubefile_default')
	if config.domain == '' {
		config_file = $tmpl('templates/peertubefile_all')
	}
	install()!
	os.mkdir_all(config.path)!

	default_html := '
	<!DOCTYPE html>
	<html>
		<head>
			<title>Peertube has now been installed.</title>
		</head>
		<body>
			Page loaded at: {{now | date "Mon Jan 2 15:04:05 MST 2006"}}
		</body>
	</html>
	'
	osal.file_write('${config.path}/index.html', default_html)!

	configuration_set(content: config_file)!
}

pub fn configuration_get() !string {
	c := osal.file_read('/etc/peertube/Peertubefile')!
	return c
}

[params]
pub struct ConfigurationArgs {
pub mut:
	content string
	path    string
	restart bool = true
}

pub fn configuration_set(args_ ConfigurationArgs) ! {
	mut args := args_
	if args.content == '' && args.path == '' {
		return error('need to specify content or path.')
	}
	if args.content.len > 0 {
		args.content = texttools.dedent(args.content)
		if !os.exists('/etc/peertube') {
			os.mkdir_all('/etc/peertube')!
		}
		osal.file_write('/etc/peertube/Peertubefile', args.content)!
	} else {
		mut p := pathlib.get_file(path: args.path, create: true)!
		content := p.read()!
		if !os.exists('/etc/peertube') {
			os.mkdir_all('/etc/peertube')!
		}
		osal.file_write('/etc/peertube/Peertubefile', content)!
	}

	if args.restart {
		restart()!
	}
}

// start peertube
pub fn start() ! {
	if !os.exists('/etc/peertube/Peertubefile') {
	}
	mut t := tmux.new()!
	mut w := t.window_new(
		name: 'peertube'
		cmd: '
			peertube run --config /etc/peertube/Peertubefile
			echo CADDY STOPPED
			/bin/bash'
	)!
}

pub fn stop() ! {
	mut t := tmux.new()!
	t.window_delete(name: 'peertube')!
	// osal.execute_silent('peertube stop') or {}
}

pub fn restart() ! {
	stop()!
	start()!
}

// if cmd_exists('peertube') {
// 	println('Peertube was already installed.')
// 	//! should we set peertube as done here !
// 	return
// }
// //TODO: better to start from a build one
// osal.execute_silent("
// 	sudo apt install -y debian-keyring debian-archive-keyring apt-transport-https gpg sudo
// 	rm -f /usr/share/keyrings/peertube-stable-archive-keyring.gpg
// 	curl -1sLfk 'https://dl.cloudsmith.io/public/peertube/stable/gpg.key' | gpg --dearmor -o /usr/share/keyrings/peertube-stable-archive-keyring.gpg
// 	curl -1sLfk 'https://dl.cloudsmith.io/public/peertube/stable/debian.deb.txt' | tee /etc/apt/sources.list.d/peertube-stable.list
// 	apt update
// 	apt install peertube
// ") or {
// 	return error('Cannot install peertube.\n${err}')
// }
