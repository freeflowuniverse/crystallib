module git3

// https://git3.com/settings/tokens
