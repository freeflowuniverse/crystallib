module docker


//https://docs.docker.com/engine/api/v1.41/#

