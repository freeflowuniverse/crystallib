module algo
