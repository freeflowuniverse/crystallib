module baobab

