module python
