module baobab
