module jobs

import freeflowuniverse.crystallib.data.params
import time
