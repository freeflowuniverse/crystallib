module openrpc_client

pub struct Animal {
	name       string
	species    string
	created_at string
}
