module models


pub struct KubernetesModel {

}

pub fn (mut km KubernetesModel)deploy(){
	println("Not Implemented")
}

pub fn (mut km KubernetesModel)delete(){
	println("Not Implemented")
}
pub fn (mut km KubernetesModel)get(){
	println("Not Implemented")
}
pub fn (mut km KubernetesModel)update(){
	println("Not Implemented")
}