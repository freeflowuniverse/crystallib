module actionsparser

// make sure that only actions are remembered linked to the actor or book and also sorted in right order
pub fn (mut actions ActionsParser) filter() ! {

}
