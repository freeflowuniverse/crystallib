module publisher

fn test_get()! {
	_ := get('')!
}