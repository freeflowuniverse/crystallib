module planner

import crystallib.texttools

// texttools.text_to_params()?
