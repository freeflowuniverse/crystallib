module rest

// todo
