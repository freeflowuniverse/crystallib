module publisher

import freeflowuniverse.crystallib.baobab.base

pub struct Collection {
	base.Base
	name string
	url string
}