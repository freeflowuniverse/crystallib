module github

//https://github.com/settings/tokens