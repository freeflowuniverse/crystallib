module main

import freeflowuniverse.crystallib.threefold.deploy 

fn main(){

}