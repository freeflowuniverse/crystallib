module gitea_client


