module bizmodel

pub struct Employee {
pub:
	name                 string
	description          string
	department           string
	cost                 string
	cost_percent_revenue f64
	nrpeople             string
	indexation           f64
	cost_center          string
	page 				 string
}


pub struct Costcenter {
pub:
	name                 string
	description          string
	department           string
}
