module blockchain

// import freeflowuniverse.crystallib.core.playbook

pub struct Controller {
}

pub fn new() !Controller {
	mut c := Controller{}
	return c
}
