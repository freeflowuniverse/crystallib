module bizmodel
