module serializers

