module planner

import freeflowuniverse.crystallib.texttools

// texttools.text_to_params()?
