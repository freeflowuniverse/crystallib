module openrpc
