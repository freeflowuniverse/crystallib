module b2

// res:=py.exec(cmd:cmd)!
