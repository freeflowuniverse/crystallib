module biz
