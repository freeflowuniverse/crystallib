module components

