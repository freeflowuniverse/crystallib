module gitea_client


struct GiteaClient {
}

