module console

import freeflowuniverse.crystallib.ui.uimodel { QuestionArgs }

pub fn (mut c UIConsole) ask_date(args QuestionArgs) string {
	panic('implement')
}

pub fn (mut c UIConsole) ask_time(args QuestionArgs) string {
	panic('implement')
}
