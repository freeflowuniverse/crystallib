module library

pub fn new() Library{
	return Library{}
}