module markdownparser

import freeflowuniverse.crystallib.core.pathlib
import freeflowuniverse.crystallib.baobab.smartid
import freeflowuniverse.crystallib.data.paramsparser

pub struct DocBase {
pub mut:
	id int //the unique id while loading of the element in the parser
	content string
	items   []DocItem [skip; str: skip]
	parent  ?DocItem [skip; str: skip]
	path    ?pathlib.Path 
	processed bool
	params ?paramsparser.Params
}

pub struct Doc {
	DocBase
pub mut:
	gid 	smartid.GID
	pre     []HtmlSource
}



[param]
pub struct HtmlSource {
pub mut:
	url         string
	path        string
	bookname    string
	chaptername string
	filename    string
	cat         HtmlSourceCat
}

enum HtmlSourceCat {
	css
	script
}


// add a css or script link to a document
//  url: is source where the data comes from, can be CDN or local link
//  path: can be relative or absolute path to the info
// 	bookname, if in memory in a book
//  chaptername, if in memory in a book
//	filename string, if in memory in a book
//  cat, is .css or .script
pub fn (mut doc Doc) pre_add(arg HtmlSource) string {
	// TODO what is this function for?
	return ''
}

type DocItem = Action | Actions | CodeBlock | Header | Html | Include | Link | Paragraph | Table | None

pub fn (mut doc Doc) wiki() string {
	mut out := ''
	for mut item in doc.items {
		match mut item {
			Table { out += item.wiki() }
			Action { out += item.wiki() }
			Actions { out += item.wiki() }
			Header { out += item.wiki() }
			Paragraph { out += item.wiki() }
			Html { out += item.wiki() }
			Include { out += item.wiki() }
			// Comment { out += item.wiki() }
			CodeBlock { out += item.wiki() }
			Link { out += item.wiki() }
			else{}
		}
	}
	return out
}

pub fn (mut doc Doc) markdown() string {
	mut out := ''
	for mut item in doc.items {
		match mut item {
			Table { out += item.wiki() }
			Action { out += item.wiki() }
			Actions { out += item.wiki() }
			Header { out += item.wiki() }
			Paragraph { out += item.markdown() }
			Html { out += item.wiki() }
			Include { out += item.wiki() }
			// Comment { out += item.wiki() }
			CodeBlock { out += item.wiki() }
			Link { out += item.markdown() }
			else{}
		}
	}
	return out
}

pub fn (mut doc Doc) html() string {
	mut out := ''
	for mut item in doc.items {
		match mut item {
			Table { out += item.html() }
			Action { out += item.html() }
			Actions { out += item.html() }
			Header { out += item.html() }
			Paragraph { out += item.html() }
			Html { out += item.html() }
			Include { out += item.html() }
			// Comment { out += item.html() }
			CodeBlock { out += item.html() }
			Link { out += item.html() }
			else{}
		}
	}
	return out
}

pub fn (mut doc Doc) save_wiki() ! {
	mut path := doc.path or {pathlib.Path{}}
	if path.path.len>0{
		path.write(doc.wiki())!
	}
}

