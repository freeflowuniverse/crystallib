module conversiontools
