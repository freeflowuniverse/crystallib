module filedb
