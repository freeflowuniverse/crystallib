module taiga
import despiegk.crystallib.crystaljson
import despiegk.crystallib.texttools
// import x.json2 { raw_decode }
import json
import time { Time }
import math { min }


enum TaskStatus { 
	//TODO: there will be many other statuses used, we have to fix, in taiga itself, make the story status as below eveywhere
	unknown
	new
	accepted
	inprogress
	verification //is called ready for test in taiga
	done
}


pub struct Task {
pub mut:
	description            string
	id                     int
	tags                   []string
	project                int
	user_story             int
	status                 TaskStatus
	assigned_to            int
	owner                  int
	created_date           Time       
	modified_date          Time        
	finished_date          Time        
	due_date               Time        
	due_date_reason        string
	subject                string
	is_closed              bool
	is_blocked             bool
	blocked_note           string
	ref                    int
	total_comments         int //TODO: why is this needed if we already have comments list? everyone can do count()?
	comments               []Comment   
	file_name              string
}

struct NewTask {
pub mut:
	subject string
	project int
}

pub fn tasks() ? {
	mut conn := connection_get()
	blocks := conn.get_json_list('tasks', '', true) ?
	println('[+] Loading $blocks.len tasks ...')
	for t in blocks {
		mut task := Task{}
		task = task_decode(t.str()) or {
			eprintln(err)
			Task{}
		}
		if task != Task{} {
			conn.task_remember(task)
		}
	}
}

// get comments in lis from task
pub fn (mut t Task) get_comments() ?[]Comment {
	t.comments = comments_get('task', t.id) ?
	return t.comments
}

pub fn task_create(subject string, project_id int) ?Task {
	mut conn := connection_get()
	task := NewTask{
		subject: subject
		project: project_id
	}
	postdata := json.encode_pretty(task)
	response := conn.post_json_str('tasks', postdata, true) ?
	mut result := task_decode(response) ?
	conn.task_remember(result)
	return result
}

pub fn task_get(id int) ?Task {
	mut conn := connection_get()
	response := conn.get_json_str('tasks/$id', '', true) ?
	mut result := task_decode(response) ?
	conn.task_remember(result)
	return result
}

pub fn task_delete(id int) ?bool {
	mut conn := connection_get()
	response := conn.delete('tasks', id) ?
	conn.task_forget(id)
	return response
}

fn task_decode(data string) ?Task {


	data_as_map := crystaljson.json_dict_any(data,false,[],[])?

	mut task:=Task{
		//TODO: put properties in		
	}

	task.comments = []


	projname:=data_as_map["project_extra_info"].as_map()["name"].str().to_upper()
	if projname.contains("ARCHIVE"){
		//this is a task linked to a project which is archived, no reason to process
		return Task{}
	}

	// println(data_as_map)

	task.created_date = parse_time(data_as_map['created_date'].str())
	task.modified_date = parse_time(data_as_map['modified_date'].str())
	task.finished_date = parse_time(data_as_map['finished_date'].str())
	task.due_date = parse_time(data_as_map['due_date'].str())
	task.file_name = texttools.name_clean(task.subject[0..min(40, task.subject.len)] + '-' + task.id.str()) + '.md'
	task.file_name = texttools.ascii_clean(task.file_name)
	if true{
		println(task.file_name)
		panic('sss')
	}	
	// task.user_story_extra_info.file_name =
	// 	texttools.name_clean(task.user_story_extra_info.subject[0..min(40, task.user_story_extra_info.subject.len)] +
	// 	'-' + task.user_story_extra_info.id.str()) + '.md'
	// task.project_extra_info.file_name =
	// 	texttools.name_clean(task.project_extra_info.slug) + '.md'
	mut conn := connection_get()
	if conn.settings.comments_task{
		task.get_comments()?
	}
	return task
}

// export template per task
pub fn (task Task) as_md(url string) string {
	mut task_md := $tmpl('./templates/task.md')
	task_md = fix_empty_lines(task_md)
	return task_md
}
