module backend

pub fn (b Backend) generate_id() string {
	return ''
}
