module markdown

pub struct Paragraph{
pub:
	content string
pub mut:
	links []Link
}

