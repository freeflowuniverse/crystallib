module openrpc

// pub struct
