module blockchain

// import freeflowuniverse.crystallib.core.actionsparser

pub struct Controller {
}

pub fn new() !Controller {
	mut c := Controller{}
	return c
}
