module play

pub fn (mut session Session) run()	! {

 	session.play_mdbook()!

}
