module openrpc

pub fn (doc OpenRPC) generate_client() {
	for method in doc.methods {
	}
}
