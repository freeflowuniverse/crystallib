module v
import freeflowuniverse.crystallib.ui.console {UIConsole}

//need to do this for each type of UI channel e.g. console, telegram, ...
type UIChannel = UIConsole

pub struct UserInteraction{
pub mut:

}