module system

[heap]
pub struct ModelFactoryBase {
pub mut:
	circle u32
	id2u32 map[string]u32
}
