module lima



