module data

//Data object for @Object
pub struct @Object {
pub mut:
	id          int
	name        string
	description string
	tags		[]string
	remarks		[]int
}