module books

pub fn new() Sites {
	return Sites{}
}
