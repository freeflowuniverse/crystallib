

module builder


// pub struct SwarmArgs{
// 	reset bool
// }

// //installs docker & swarm
// fn (mut node Node) ubuntu_update(args SwarmArgs) ?{

// 	cmd := '
// 		set -ex
// 		apt update
// 		apt upgrade -y
// 		apt autoremove -y
// 		'

// 	node.exec({cmd:cmd,cache:3600*12})?

// }
