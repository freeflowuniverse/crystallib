module tfrobot

fn test_new() {
	bot := new()!
}
