
module actors
