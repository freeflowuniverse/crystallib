module doctreemodel

pub struct ObjNotFound {
	Error
pub:
	pointer Pointer
}

