module jobs

import freeflowuniverse.crystallib.params { Params }
import time
