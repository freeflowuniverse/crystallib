module library

import freeflowuniverse.crystallib.books.chapters


[heap]
pub struct Library {
pub mut:
	chapters  []chapters.Chapter
}

