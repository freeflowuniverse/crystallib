module postgresql

// import freeflowuniverse.crystallib.osal
// import freeflowuniverse.crystallib.ui.console
// import freeflowuniverse.crystallib.installers.virt.docker

// pub fn requirements() ! {
// 	if !osal.done_exists('postgres_install') {
// 		panic('to implement, check is ubuntu and then install, for now only ubuntu')
// 		osal.package_install('libpq-dev,postgresql-client')!
// 		osal.done_set('postgres_install', 'OK')!
// 		console.print_header('postgresql installed')
// 	} else {
// 		console.print_header('postgresql already installed')
// 	}
// }
