

module main

fn do() ! {



}

fn main() {
	do() or { panic(err) }
}
