module main

pub fn testfunction(param string) string {
	return param
}
