module core
