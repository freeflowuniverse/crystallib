module jsonschema
