module base

pub struct Base {
pub mut:
	id u32
}
