module code


// const actor_name = 'testactor'
// const actor_path = '${os.dir(@FILE)}/testdata/${actor_name}'

const testactor := Actor{}

pub fn test_write() ! {
	// testactor.write('')!
}