module main

import freeflowuniverse.crystallib.keysafe.secp256k1

fn main() {
	println("Coucou")
}
