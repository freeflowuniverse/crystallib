module testtools

struct TestRun {
}
