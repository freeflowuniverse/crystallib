module griddriver

pub struct Client {
	mnemonic  string
	substrate string
	relay     string
}

// TODO: add the rest of griddriver functionalities
