module couchdb


//see http://127.0.0.1:5984/_utils/docs/intro/api.html#replication


pub fn (mut cl CouchDBInstance) replication_get(...)!{

}

pub fn (mut cl CouchDBInstance) replication_add(...)!{

}

pub fn (mut cl CouchDBInstance) replication_delete(...)!{

}

pub fn (mut cl CouchDBInstance) replication_list(...)!{

}
