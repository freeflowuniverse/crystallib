module main

// method_with_description shows that the parser can parse a method's description
// from its comments, even if the comments are multiline.
pub fn method_with_description(name string) {}
