module investorsimulator

pub struct CapTable{
	
}