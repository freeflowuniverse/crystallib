module backoffice

// import freeflowuniverse.protocolme.organization
// import freeflowuniverse.crystallib.core.texttools

// TODO circle_add

// TODO circle_end
/*
// Find a specific Group
pub fn (mut memdb MemDB) circle_find(circle_name string) ?&organization.Group {
	shortname := texttools.name_fix_no_underscore_no_ext(circle_name)

	if shortname in data.circles {
		return data.circles[shortname]
	}
	return error('Could not find circle with name: $shortname')
}
*/
