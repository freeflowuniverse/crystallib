module books
