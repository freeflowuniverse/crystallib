module schedule

import freeflowuniverse.crystallib.baobab.base

// pub struct Event {
// 	base.Base
// pub mut:
// 	event_name string
// }