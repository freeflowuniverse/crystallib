module data

//Data object for Story
pub struct Story {
pub mut:
	id          int
	name        string
	description string
	tags		[]string
	remarks		[]int
}