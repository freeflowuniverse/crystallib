module imagemagick

fn install() ? {
	if !installed() {
		cmd := 'brew install imagemagick'
	}
}
