module taiga

//all internal

// fn (mut h TaigaConnection) user_get(id int)? &User{

// }

// fn (mut h TaigaConnection) project_get(id int)? &Project{

// }

// fn (mut h TaigaConnection) story_get(id int)? &Story{

// }

// fn (mut h TaigaConnection) epic_get(id int)? &Epic{

// }

// fn (mut h TaigaConnection) task_get(id int)? &Task{

// }


// fn (mut h TaigaConnection) user_remember(obj User){
// 	//check obj exists in connection, if yes, update & return
// 	//make sure to remeber the reference !!!

// }

// //TODO: do same for other objects