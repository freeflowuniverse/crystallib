module ourserver

const (
	tcp_server_port = 2223
)
