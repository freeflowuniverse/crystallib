module backoffice


