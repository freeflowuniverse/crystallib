module archiver

struct FList {
}

struct FListDir {
	nr   u32
	name string
}

struct FListFile {
	nr   u32
	name string
}
