module heroencoder
