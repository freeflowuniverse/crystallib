
module tfgrid3deployer

import json
import freeflowuniverse.crystallib.data.encoder


pub struct WebName {
pub mut:
	name        string

}
