module griddriver

pub struct Client {
	substrate string
	mnemonic  string
	relay     string
}

// TODO: add the rest of griddriver functionalities
