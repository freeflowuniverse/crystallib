module books

pub fn new() Sites {
	mut sites := Sites{}
	sites.config = Config{}
	return sites
}
