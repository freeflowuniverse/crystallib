module auth

// fn get_session(mut ctx vweb.Context) bool {
// 	// impelement your own logic to get the user

// 	refresh_token := app.get_cookie('token') or { '' }

// 	user := User{
// 		session_id: '123456'
// 		name: 'Vweb'
// 	}

// 	// set the user
// 	ctx.set_value('user', user)
// 	return true
// }
