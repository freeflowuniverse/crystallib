module crypt
