module collection

import freeflowuniverse.crystallib.core.pathlib { Path }
import freeflowuniverse.crystallib.data.doctree3.collection.data
import freeflowuniverse.crystallib.core.texttools

@[heap]
pub struct Collection {
pub:
	name string @[required]
pub mut:
	path   Path                  @[required]
	pages  map[string]&data.Page
	files  map[string]&data.File
	images map[string]&data.File
	errors []CollectionError
	heal   bool = true
}

@[params]
pub struct CollectionNewArgs {
mut:
	name string @[required]
	path string @[required]
	heal bool = true // healing means we fix images, if selected will automatically load, remove stale links
	load bool = true
}

// get a new collection
pub fn new(args_ CollectionNewArgs) !Collection {
	mut args := args_
	args.name = texttools.name_fix(args.name)

	mut pp := pathlib.get_dir(path: args.path)! // will raise error if path doesn't exist
	mut collection := Collection{
		name: args.name
		path: pp
		heal: args.heal
	}

	if args.load {
		collection.scan()!
	}

	return collection
}
