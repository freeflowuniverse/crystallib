module main

import despiegk.crystallib.vredis2

fn main() {
	vredis2.redis_encode_test()
}
