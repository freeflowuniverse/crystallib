
module components
import db.sqlite
import nedpals.vex.ctx
import freeflowuniverse.crystallib.core.texttools

pub fn html_pre(req &ctx.Req)!string{
	out:='
	<!DOCTYPE html>
	<html lang="en">
	<head>
		<meta charset="UTF-8">
		<meta name="viewport" content="width=device-width, initial-scale=1.0">
		<title>Sample Form</title>
		<script src="https://cdn.tailwindcss.com"></script>
	</head>
	<body>
	'
	return texttools.dedent(out)

}

pub fn html_post(req &ctx.Req)!string{
	out:='
	</body>
	</html>
	'
	return texttools.dedent(out)
}



