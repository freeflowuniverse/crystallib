module people


pub struct Country { 
pub mut:
	name  		string
	codes 		[]string
}


