module actionsparser

import os

fn test_filter() {

}

