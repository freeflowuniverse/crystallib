module main

import regex {RE,regex_opt}

pub struct EmptyRegex {
}

type OurRegex = RE | EmptyRegex

pub struct ListArgs {
pub mut:
	regex	  OurRegex
}


fn main(){

	query := r'(c(pa)+z ?)+'
	mut re := regex_opt(query) or { panic(err) }

	item := "sss"
	mut la := ListArgs{
		regex:re
	}

	mut r:=la.regex
	if r is RE{
		println(r)
		println(r.matches_string(item))
	}

    // match r {
    //     RE { r.matches_string(item) }
    //     else {}
    // }	

}
