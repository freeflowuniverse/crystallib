module zerohub

const secret="6Pz6giOpHSaA3KdYI6LLpGSLmDmzmRkVdwvc7S-E5PVB0-iRfgDKW9Rb_ZTlj-xEW4_uSCa5VsyoRsML7DunA1sia3Jpc3RvZi4zYm90IiwgMTY3OTIxNTc3MF0="

fn test_main() ? {

	mut cl := new(secret:secret)!

	// flists := cl.get_flists()!
	// println(flists)

	// repos := cl.get_repos()!
	// println(repos)

	// files := cl.get_files()!
	// println(files)

	// flists := cl.get_repo_flists('omarabdulaziz.3bot')!
	// println(flists)

	// flist_data := cl.get_flist_dump('omarabdulaziz.3bot', 'omarabdul3ziz-obuntu-zinit.flist')!
	// println(flist_data)

}