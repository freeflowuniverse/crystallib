module gittools

import os
import freeflowuniverse.crystallib.osal.sshagent
import freeflowuniverse.crystallib.core.texttools
import freeflowuniverse.crystallib.core.pathlib

fn test_check() {
}

fn test_addr_from_path() {
}

fn test_path() {
}

fn test_path_account() {
}

fn test_url_get() {
}

fn test_url_ssh_get() {
}

fn test_url_http_get() {
}

fn test_url_http_with_branch_get() {
}

fn test_str() {
}
