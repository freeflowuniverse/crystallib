module main
import freeflowuniverse.crystallib.builder
import installers.mdbook
import installers.caddy

fn do() ? {
	// shortcut to install the base
	mut builder := builder.new()
	mut node := builder.node_new(ipaddr:"185.206.122.153",name:"kds")?
	caddy.get_install(mut node)?
	mdbook.get_install(mut node)?
}

fn main() {
	do() or { panic(err) }
}
