module library

