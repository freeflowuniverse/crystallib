module twinsafe

//TODO: create 3 tables, one for othertwin, one for mytwin, one for myconfig