module elements

import freeflowuniverse.crystallib.core.smartid

@[heap]
pub struct Doc {
	DocBase
pub mut:
	gid smartid.GID
	pre []HtmlSource
}

// add a css or script link to a document
//  url: is source where the data comes from, can be CDN or local link
//  path: can be relative or absolute path to the info
// 	bookname, if in memory in a book
//  chaptername, if in memory in a book
//	filename string, if in memory in a book
//  cat, is .css or .script
pub fn (mut self Doc) pre_add(arg HtmlSource) string {
	return ''
}

@[param]
pub struct HtmlSource {
pub mut:
	url         string
	path        string
	bookname    string
	chaptername string
	filename    string
	cat         HtmlSourceCat
}

enum HtmlSourceCat {
	css
	script
}

@[params]
pub struct DocNewArgs {
pub mut:
	gid     smartid.GID
	pre     []HtmlSource
	content string
}

pub fn doc_new(args DocNewArgs) !Doc {
	mut d := Doc{
		gid: args.gid
		pre: args.pre
	}
	return d
}

pub fn (mut self Doc) remove_empty_elements() ! {
	mut to_delete := []int{}
	for id, element in self.children {
		// remove the elements which are empty
		if element.content.trim_space() == '' {
			to_delete << id
		}
	}

	self.delete_from_children(to_delete)
}
