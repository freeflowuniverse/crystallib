module serializers
