module installers
