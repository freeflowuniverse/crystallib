module couchdb

// see http://127.0.0.1:5984/_utils/docs/intro/api.html#documents attachments

// make sure we return as binary

// QUESTION: how should we deal with big documents

pub fn (mut cl CouchDBInstance) attachment_get() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) attachment_add() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) attachment_delete() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) attachment_list() ! {
	panic('implement')
}
