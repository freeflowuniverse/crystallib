module zola

fn test_section_export() {
	section := Section{}
	section.export('test')!
<<<<<<< HEAD
}
=======
}
>>>>>>> e61681d (example fix wip)
