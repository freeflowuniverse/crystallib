module encoder
