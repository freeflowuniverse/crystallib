module sshagent

// fn listsplit(key string) string {
// 	if key.trim(' ') == '' {
// 		return ''
// 	}
// 	if key.contains(' ') {
// 		splitted := key.split(' ')
// 		return splitted[splitted.len].replace('.pub', '')
// 	}
// 	return key
// }
