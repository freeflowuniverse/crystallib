module msgbus
