module clients
