module sshagent


// [params]
// pub struct KeyExistsArgs{
// 	pubkey string
// 	privkey string
// 	pubkey_path string
// 	privkey_path string
// 	name string
// }

// pub fn key_exists(args) KeyExistsArgs) bool {
// 	pubkeys:=pubkeys_get()
// 	return pubkey in pubkeys
// }

//TODO: kristof refactor sshagent