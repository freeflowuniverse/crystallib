module secp256k1

#include "@VMODROOT/secp256k1.h"

#flag @VMODROOT/secp256k1.o
#flag -lsecp256k1

fn main() {
	println("Hello World")
}
