module petstore_client

struct Pet {
	name string
	tag string
	id int
}