module tfgrid

// see https://github.com/threefoldtech/zos/tree/provision-engine-cleanup/pkg/gridtypes
