module vdc

pub struct VM {
pub mut:
	name        string
	description string
	vms         []DISK
}
