module blockchain

// import freeflowuniverse.crystallib.baobab.actions


pub struct Controller {
}

pub fn new() !Controller {
	mut c:=Controller{}
	return c
}

