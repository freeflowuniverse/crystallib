module components