module knowledgetree

pub fn new() Tree {
	return Tree{}
}
