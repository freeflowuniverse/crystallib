module osal

fn test_new_osal() {
	o := new()!
}