module planner

import despiegk.crystallib.texttools

// texttools.text_to_params()?
