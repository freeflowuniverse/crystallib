module bizmodel

pub struct BizModelArgs{
pub mut:
	name string
	data_path string
}