module couchdb

// see http://127.0.0.1:5984/_utils/docs/intro/api.html#replication

pub fn (mut cl CouchDBInstance) replication_get() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) replication_add() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) replication_delete() ! {
	panic('implement')
}

pub fn (mut cl CouchDBInstance) replication_list() ! {
	panic('implement')
}
