
module tfgrid3deployer

import json
import freeflowuniverse.crystallib.data.encoder


pub struct ZDB {
pub mut:
	name        string
}

