module filedb

