module docker
import freeflowuniverse.crystallib.params {Params}

[params]
pub struct BuildArgs{
pub mut:
	args Params
	reset bool
	strict bool
}
