module downloader

// pub fn url_is_git_repo(url string) bool {

// 	// url is Git Transport Protocol
// 	// git://host.xz/path/to/repo.git/ or git://host.xz/~user/path/to/repo.git/
// 	if url.starts_with('git://') {
// 		if url.trim_string_left('git://').count('/') < 2 {
// 			return false
// 		}
// 		// TODO: perform more checks
// 		return true
// 	}

// 	http_schema := url.starts_with('http://') || u.starts_with('https://')

// }
