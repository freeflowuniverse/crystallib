module macros

import time
import freeflowuniverse.crystallib.core.texttools

fn macro_time(mut state LineProcessorState, mut macro texttools.MacroObj) ? {
	mut out := []string{}

	now := time.now()
	out << 'Generated on `' + now.format_ss() + '`'

	state.lines_server << out
}
