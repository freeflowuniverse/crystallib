module hero

import freeflowuniverse.crystallib.baobab.actions

// recursive include of actions
fn (mut s Session) actions_git(myactions []actions.Action) ! {
}
