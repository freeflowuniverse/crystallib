module penapp

fn pen_run(){

}