module rest


const version = "1"
