module installers

// TODO: how to deal with environment os.env
