module keydb

// make BUILD_TLS=no ENABLE_FLASH=yes  V=1
// export LDFLAGS="-L/opt/homebrew/opt/openssl@3/lib -L/opt/homebrew/opt/zstd"
// export CPPFLAGS="-I/opt/homebrew/opt/openssl@3/include -I/opt/homebrew/opt/zstd/include"
// https://github.com/Snapchat/KeyDB

// https://github.com/Snapchat/ModJS
