module sendGrid

import net.http