module pen

fn pen_run(){

}