module console

pub fn clear(){
	print("\033[2J")
}