module publisher_config

// // {
// //   "name": "incachain",
// //   "cat": 0,
// //   "descr": "",
// //   "depends": []
// // }
// pub struct SiteConfigLocal {
// pub mut:
// 	name       string
// 	cat        SiteCat
// 	descr      string
// 	depends []SiteDependency
// }



// pub struct SiteDependency {
// pub mut:
// 	url       string
// 	path        string  //path in the git repo as defined by the url
// 	fs_path	  string    //path as on fs, can be local to the location of this config file
// 	branch      string
// }



