module pmdb

import freeflowuniverse.protocolme.models.people
import freeflowuniverse.protocolme.models.system
// import freeflowuniverse.protocolme.models.backoffice.organization
import time



[heap]
pub struct MemDB {
pub mut:
	
}


pub fn new() MemDB {
	return MemDB{}
}
